// ID
module Shift_Left_Two_32(
    data_i,
    data_o
    );

// TO DO
  
     
endmodule
