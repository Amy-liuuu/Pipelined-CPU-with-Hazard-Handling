// ID
module MUX_2to1(
               data0_i,
               data1_i,
               select_i,
               data_o
               );

// TO DO


endmodule      
